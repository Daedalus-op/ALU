module multiplier (
  input  [1:0] a, b,
  output [3:0]product
);
  wire p[3:0], q[3:0];
  reg sum[3:0];

endmodule
