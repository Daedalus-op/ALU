module alu_tb;
  
reg clk;
wire y;

endmodule
